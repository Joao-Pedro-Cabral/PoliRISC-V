
package macros_pkg;
  `default_nettype none
  timeunit 1ns / 1ns;
endpackage
