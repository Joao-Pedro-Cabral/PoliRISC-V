../../simulation/board.vh