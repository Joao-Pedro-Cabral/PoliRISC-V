
package macros_pkg;
  timeunit 1ns / 1ns;
endpackage
