`define LITEX_
