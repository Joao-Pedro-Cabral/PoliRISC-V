
module Dataflow_tb();

endmodule