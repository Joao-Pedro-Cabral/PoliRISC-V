`define ZICSR 
`define TrapReturn 
