../../../simulation/macros.vh