`define UART_0 
