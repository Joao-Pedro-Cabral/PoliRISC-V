`define UART_0
