import hazard_unit_pkg::*;
import dataflow_pkg::*;

module dataflow #(
    parameter integer DATA_SIZE = 32
) (
    // Common
    input wire clock,
    input wire reset,
    // Instruction Memory
    input wire [DATA_SIZE-1:0] inst,
    output wire [DATA_SIZE-1:0] inst_mem_addr,
    // Data Memory
    input wire [DATA_SIZE-1:0] rd_data,
    output wire [DATA_SIZE-1:0] wr_data,
    output wire [DATA_SIZE-1:0] data_mem_addr,
    // From Memory Unit
    input logic mem_busy,
    // From Control Unit
    input wire alua_src,
    input wire alub_src,
`ifdef RV64I
    input wire aluy_src,
`endif
    input wire [3:0] alu_src,
    input wire sub,
    input wire arithmetic,
    input wire alupc_src,
    input wire pc_src,
    input wire pc_en,
    input wire [1:0] wr_reg_src,
    input wire wr_reg_en,
    input wire ir_en,
    input wire mem_addr_src,
    input forwarding_type_t forwarding_type,
    // Interrupts/Exceptions from UC
    input wire ecall,
    input wire illegal_instruction,
    // Trap Return
    input wire mret,
    input wire sret,
    // Interrupts from Memory
    input wire external_interrupt,
    input wire [DATA_SIZE-1:0] mem_msip,
    input wire [63:0] mem_mtime,
    input wire [63:0] mem_mtimecmp,
    input wire csr_wr_en,
    input wire [1:0] csr_op,
    input wire csr_imm,
    // To Control Unit
    output wire [6:0] opcode,
    output wire [2:0] funct3,
    output wire [6:0] funct7,
    output wire zero,
    output wire negative,
    output wire carry_out,
    output wire overflow,
    output wire csr_addr_exception,
    output wire [1:0] privilege_mode,
    // From Forwarding Unit
    input forwarding_t forward_rs1_id,
    input forwarding_t forward_rs2_id,
    input forwarding_t forward_rs1_ex,
    input forwarding_t forward_rs2_ex,
    input forwarding_t forward_rs2_mem,
    // To Forwarding Unit
    output forwarding_type_t forwarding_type_id,
    output forwarding_type_t forwarding_type_ex,
    output forwarding_type_t forwarding_type_mem,
    output logic reg_we_mem,
    output logic reg_we_wb,
    output logic zicsr_ex,
    output logic [4:0] rd_ex,
    output logic [4:0] rd_mem,
    output logic [4:0] rd_wb,
    output logic [4:0] rs1_id,
    output logic [4:0] rs2_id,
    output logic [4:0] rs1_ex,
    output logic [4:0] rs2_ex,
    output logic [4:0] rs2_mem,
    // From Hazard Unit
    input logic stall_if,
    input logic stall_id,
    input logic flush_id,
    input logic flush_ex,
    // To Hazard Unit
    output hazard_t hazard_type,
    output rs_used_t rs_used,
    output logic [4:0] rs1_id,
    output logic [4:0] rs2_id,
    output logic [4:0] rd_ex,
    output logic [4:0] rd_mem,
    output logic reg_we_ex,
    output logic reg_we_mem,
    output logic mem_rd_en_ex,
    output logic mem_rd_en_mem,
    output logic zicsr_ex,
    output logic store_id
);

  // Pipeline registers
  if_id_t                  if_id_reg;
  id_ex_t                  id_ex_reg;
  ex_mem_t                 ex_mem_reg;
  mem_wb_t                 mem_wb_reg;

  // Fios intermediários
  // Register File
  wire     [          4:0] rs1_addr;
  wire     [DATA_SIZE-1:0] rs1;
  wire     [DATA_SIZE-1:0] rs2;
  wire     [DATA_SIZE-1:0] rd;
  // Extensor de Imediato
  wire     [DATA_SIZE-1:0] immediate;
  // ULA
  wire     [DATA_SIZE-1:0] aluA;
  wire     [DATA_SIZE-1:0] aluB;
  wire     [DATA_SIZE-1:0] aluY;
  wire     [DATA_SIZE-1:0] muxaluY_out;  // aluY or sign_extended(aluY[31:0])
  // Somador PC + 4
  wire     [DATA_SIZE-1:0] pc_plus_4;
  wire     [DATA_SIZE-1:0] cte_4 = 4;
  // Somador PC + Imediato
  wire     [DATA_SIZE-1:0] pc_plus_immediate;
  // PC
  wire     [DATA_SIZE-1:0] pc;
  reg      [DATA_SIZE-1:0] new_pc;
  // Instruction Register(IR)
  wire     [         31:0] ir;
  // CSR
  wire     [DATA_SIZE-1:0] trap_addr;
  wire                     _trap;
  wire     [          1:0] _privilege_mode;
  // Trap Return
  wire     [DATA_SIZE-1:0] mepc;
  wire     [DATA_SIZE-1:0] sepc;
  // ZICSR
  wire     [DATA_SIZE-1:0] csr_rd_data;
  wire     [DATA_SIZE-1:0] csr_mask_rd_data;
  wire     [DATA_SIZE-1:0] csr_wr_data;
  wire     [DATA_SIZE-1:0] csr_aux_wr;

  // IF stage
  always_ff @(posedge clock iff (~stall_if && ~mem_busy) or posedge reset) begin
    if (reset) if_id_reg <= '0;
    else if (flush_id) if_id_reg <= '0;
    else begin
      if_id_reg.pc <= new_pc;
      if_id_reg.pc_plus_4 <= pc_plus_4;
      if_id_reg.inst <= inst;
    end
  end

  always_comb begin
    if (_trap) new_pc = trap_addr;
    else if (mret) new_pc = mepc;
    else if (sret) new_pc = sepc;
    else if (pc_src) new_pc = pc_plus_immediate;
    else new_pc = pc_plus_4;
  end

  // PC
  register_d #(
      .N(DATA_SIZE),
      .reset_value(0)
  ) pc_register (
      .clock(clock),
      .reset(reset),
      .enable(~stall_if && ~mem_busy),
      .D(new_pc),
      .Q(pc)
  );

  // Memory
  assign inst_mem_addr = pc;
  // IF stage

  // Instanciação de Componentes
  // Register File
  gen_mux #(
      .size(DATA_SIZE),
      .N(2)
  ) mux11 (
      .A({pc_plus_4, rd_data, csr_mask_rd_data, muxaluY_out}),
      .S(wr_reg_src),
      .Y(rd)
  );
  // caso seja realizada uma leitura do SEIP(9) é preciso realizar o OR com o external_interrupt
  assign csr_mask_rd_data[8:0] = csr_rd_data[8:0];
  assign csr_mask_rd_data[9] = (ir[31:20] == 12'h344 || ir[31:20] == 12'h144)
                                            ? (csr_rd_data[9] | external_interrupt)
                                            : csr_rd_data[9];
  assign csr_mask_rd_data[DATA_SIZE-1:10] = csr_rd_data[DATA_SIZE-1:10];

  register_file #(
      .size(DATA_SIZE),
      .N(5)
  ) int_reg_state (
      .clock(clock),
      .reset(reset),
      // You can't write an illegal value coming from CSR
      .write_enable(wr_reg_en && !(wr_reg_src == 2'b01 && csr_addr_exception)),
      .read_address1(rs1_addr),
      .read_address2(ir[24:20]),
      .write_address(ir[11:7]),
      .write_data(rd),
      .read_data1(rs1),
      .read_data2(rs2)
  );
  // ULA
`ifdef RV64I
  assign aluA = alua_src ? pc : (aluy_src ? {{32{rs1[31]}}, rs1[31:0]} : rs1);
  assign aluB = alub_src ? immediate : (aluy_src ? {{32{rs2[31]}}, rs2[31:0]} : rs2);
  assign muxaluY_out[DATA_SIZE-1:32] = aluy_src ? {32{aluY[31]}} : aluY[DATA_SIZE-1:32];
`else
  assign aluA = alua_src ? pc : rs1;
  assign aluB = alub_src ? immediate : rs2;
`endif

  ULA #(
      .N(DATA_SIZE)
  ) alu (
      .A(aluA),
      .B(aluB),
      .seletor(alu_src),
      .sub(sub),
      .arithmetic(arithmetic),
      .Y(aluY),
      .zero(zero),
      .negative(negative),
      .carry_out(carry_out),
      .overflow(overflow)
  );
  // Somador PC + 4
  sklansky_adder #(
      .INPUT_SIZE(DATA_SIZE)
  ) pc_4 (
      .A(pc),
      .B(cte_4),
      .c_in(1'b0),
      .c_out(),
      .S(pc_plus_4)
  );
  // Somador PC + Imediato
  sklansky_adder #(
      .INPUT_SIZE(DATA_SIZE)
  ) pc_immediate (
      .A(alupc_src ? {rs1[DATA_SIZE-1:1], 1'b0} : pc),
      .B({immediate[DATA_SIZE-1:1], 1'b0}),
      .c_in(1'b0),
      .c_out(),
      .S(pc_plus_immediate)
  );
  // Immediate Extender
  immediate_extender #(
      .N(DATA_SIZE)
  ) estende_imediato (
      .instruction(ir),
      .immediate  (immediate)
  );
  // Instruction Register -> Borda de Descida!
  register_d #(
      .N(32),
      .reset_value(0)
  ) instru_register (
      .clock(clock),
      .reset(reset),
      .enable(ir_en),
      .D(rd_data[31:0]),
      .Q(ir)
  );
  // CSR
  CSR csr_bank (
      .clock(clock),
      .reset(reset),
      .trap_en(~stall_if && ~mem_busy),
      // Interrupt/Exception Signals
      .ecall(ecall),
      .illegal_instruction(illegal_instruction),
      .external_interrupt(external_interrupt),
      .mem_msip(|mem_msip),
      .mem_mtime(mem_mtime),
      .mem_mtimecmp(mem_mtimecmp),
      .trap_addr(trap_addr),
      .trap(_trap),
      .privilege_mode(_privilege_mode),
      .addr_exception(csr_addr_exception),
      .pc(pc),
      .instruction(ir),
      // CSR RW interface
      .wr_en(csr_wr_en & (~csr_op[1] | (|ir[19:15]))),
      .addr(ir[31:20]),
      .wr_data(csr_wr_data),
      .rd_data(csr_rd_data),
      // TrapReturn
      .mret(mret),
      .sret(sret),
      .mepc(mepc),
      .sepc(sepc)
  );


  // Atribuições intermediárias
  // Mascarar LUI no Rs1
  assign rs1_addr = ir[19:15] & {5{(~(ir[4] & ir[2]))}};
  assign muxaluY_out[31:0] = aluY[31:0];

  // Zicsr
  assign csr_aux_wr = csr_imm ? $unsigned(ir[19:15]) : rs1;
  assign csr_wr_data = csr_op[1] ? (csr_op[0] ? (csr_rd_data & (~csr_aux_wr))
                        : (csr_rd_data | csr_aux_wr)) : csr_aux_wr;

  // Saídas
  // Memory
  assign wr_data = rs2;
  // Control Unit
  assign opcode = ir[6:0];
  assign funct3 = ir[14:12];
  assign funct7 = ir[31:25];
  assign privilege_mode = _privilege_mode;

endmodule
