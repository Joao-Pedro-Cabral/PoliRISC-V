../../simulation/extensions.vh