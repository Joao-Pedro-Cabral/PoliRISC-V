`define RV64I
