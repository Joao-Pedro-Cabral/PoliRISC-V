`define TrapReturn
`define M
`define ZICSR
