/home/joao/Documents/Poli/IC/RISC-V/2023s1-sd2-risc-v/simulation/macros.vh